//DESIGN "test1"
//DATE "Tue Oct 31 10:32:34 2023"
//VENDOR "NanoXplore"
//PROGRAM "Impulse"
//VERSION "v23.3.0.2"

module test1 (
  input          i_A,
  input  [7:0]   i_data,
  output [7:0]   o_data,
  output [7:0]   o_data1
);

wire data1_0;
wire data1_1;
wire data1_2;
wire data1_3;
wire data1_4;
wire data1_5;
wire data1_6;
wire data1_7;
wire data_0;
wire data_1;
wire data_2;
wire data_3;
wire data_4;
wire data_5;
wire data_6;
wire data_7;
wire r_i_A;
wire r_i_data_0;
wire r_i_data_1;
wire r_i_data_2;
wire r_i_data_3;
wire r_i_data_4;
wire r_i_data_5;
wire r_i_data_6;
wire r_i_data_7;


NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1110010011100100)
  )
  i_LOGIC_lut_10 (
   .I1(r_i_A)
  ,.I2(data_2)
  ,.I3(r_i_data_2)
  ,.I4(1'b0)
  ,.O(data_2)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1101100011011000)
  )
  i_LOGIC_lut_6 (
   .I1(r_i_A)
  ,.I2(data1_6)
  ,.I3(r_i_data_6)
  ,.I4(1'b0)
  ,.O(data1_6)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1101110110001000)
  )
  i_LOGIC_lut_11 (
   .I1(r_i_A)
  ,.I2(r_i_data_3)
  ,.I3(1'b0)
  ,.I4(data_3)
  ,.O(data_3)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111000011001100)
  )
  i_LOGIC_lut_13 (
   .I1(1'b0)
  ,.I2(data_5)
  ,.I3(r_i_data_5)
  ,.I4(r_i_A)
  ,.O(data_5)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111101001010000)
  )
  i_LOGIC_lut_2 (
   .I1(r_i_A)
  ,.I2(1'b0)
  ,.I3(r_i_data_2)
  ,.I4(data1_2)
  ,.O(data1_2)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111000011001100)
  )
  i_LOGIC_lut_15 (
   .I1(1'b0)
  ,.I2(data_7)
  ,.I3(r_i_data_7)
  ,.I4(r_i_A)
  ,.O(data_7)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111010110100000)
  )
  i_LOGIC_lut_8 (
   .I1(r_i_A)
  ,.I2(1'b0)
  ,.I3(r_i_data_0)
  ,.I4(data_0)
  ,.O(data_0)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111110000110000)
  )
  i_LOGIC_lut_9 (
   .I1(1'b0)
  ,.I2(r_i_A)
  ,.I3(data_1)
  ,.I4(r_i_data_1)
  ,.O(data_1)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1111010110100000)
  )
  i_LOGIC_lut_14 (
   .I1(r_i_A)
  ,.I2(1'b0)
  ,.I3(r_i_data_6)
  ,.I4(data_6)
  ,.O(data_6)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1101100011011000)
  )
  i_LOGIC_lut_0 (
   .I1(r_i_A)
  ,.I2(data1_0)
  ,.I3(r_i_data_0)
  ,.I4(1'b0)
  ,.O(data1_0)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1110010011100100)
  )
  i_LOGIC_lut_3 (
   .I1(r_i_A)
  ,.I2(r_i_data_3)
  ,.I3(data1_3)
  ,.I4(1'b0)
  ,.O(data1_3)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1011101110001000)
  )
  i_LOGIC_lut_1 (
   .I1(data1_1)
  ,.I2(r_i_A)
  ,.I3(1'b0)
  ,.I4(r_i_data_1)
  ,.O(data1_1)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1101100011011000)
  )
  i_LOGIC_lut_12 (
   .I1(r_i_A)
  ,.I2(r_i_data_4)
  ,.I3(data_4)
  ,.I4(1'b0)
  ,.O(data_4)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1010101011110000)
  )
  i_LOGIC_lut_5 (
   .I1(data1_5)
  ,.I2(1'b0)
  ,.I3(r_i_data_5)
  ,.I4(r_i_A)
  ,.O(data1_5)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1110010011100100)
  )
  i_LOGIC_lut_4 (
   .I1(r_i_A)
  ,.I2(r_i_data_4)
  ,.I3(data1_4)
  ,.I4(1'b0)
  ,.O(data1_4)
);

NX_LUT
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  #(
   .lut_table(16'b1010101011110000)
  )
  i_LOGIC_lut_7 (
   .I1(data1_7)
  ,.I2(1'b0)
  ,.I3(r_i_data_7)
  ,.I4(r_i_A)
  ,.O(data1_7)
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[0]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB9_D10P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_0_iob (
   .O(r_i_data_0)
  ,.C(1'b0)
  ,.IO(i_data[0])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[2]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB7_D14")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_2_iob (
   .O(r_i_data_2)
  ,.C(1'b0)
  ,.IO(i_data[2])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[6]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB1_D06")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_6_iob (
   .O(r_i_data_6)
  ,.C(1'b0)
  ,.IO(i_data[6])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[1]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB3_D15N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_1_iob (
   .O(r_i_data_1)
  ,.C(1'b0)
  ,.IO(i_data[1])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_A")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB4_D03P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_A_iob (
   .O(r_i_A)
  ,.C(1'b0)
  ,.IO(i_A)
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[5]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB10_D15N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_5_iob (
   .O(r_i_data_5)
  ,.C(1'b0)
  ,.IO(i_data[5])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[3]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB2_D14P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_3_iob (
   .O(r_i_data_3)
  ,.C(1'b0)
  ,.IO(i_data[3])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[4]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB5_D08P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_4_iob (
   .O(r_i_data_4)
  ,.C(1'b0)
  ,.IO(i_data[4])
);

NX_IOB_I
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£i_data[7]")
  // alias_vhdl("NX_IOB_I")
  // alias_vlog("")
  #(
   .location("IOB3_D09P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d1)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_i_data_7_iob (
   .O(r_i_data_7)
  ,.C(1'b0)
  ,.IO(i_data[7])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[5]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB11_D13P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_5_iob (
   .I(data1_5)
  ,.C(1'b1)
  ,.IO(o_data1[5])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[3]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB13_D10N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_3_iob (
   .I(data_3)
  ,.C(1'b1)
  ,.IO(o_data[3])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[3]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB2_D13N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_3_iob (
   .I(data1_3)
  ,.C(1'b1)
  ,.IO(o_data1[3])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[0]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB3_D13N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_0_iob (
   .I(data1_0)
  ,.C(1'b1)
  ,.IO(o_data1[0])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[1]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB9_D04P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_1_iob (
   .I(data1_1)
  ,.C(1'b1)
  ,.IO(o_data1[1])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[7]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB13_D02N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_7_iob (
   .I(data1_7)
  ,.C(1'b1)
  ,.IO(o_data1[7])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[6]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB8_D02N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_6_iob (
   .I(data1_6)
  ,.C(1'b1)
  ,.IO(o_data1[6])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[2]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB8_D16N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_2_iob (
   .I(data1_2)
  ,.C(1'b1)
  ,.IO(o_data1[2])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[7]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB10_D00P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_7_iob (
   .I(data_7)
  ,.C(1'b1)
  ,.IO(o_data[7])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[4]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB3_D00N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_4_iob (
   .I(data_4)
  ,.C(1'b1)
  ,.IO(o_data[4])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[6]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB2_D06P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_6_iob (
   .I(data_6)
  ,.C(1'b1)
  ,.IO(o_data[6])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[1]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB3_D14N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_1_iob (
   .I(data_1)
  ,.C(1'b1)
  ,.IO(o_data[1])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[5]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB2_D16N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_5_iob (
   .I(data_5)
  ,.C(1'b1)
  ,.IO(o_data[5])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[0]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB0_D05")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_0_iob (
   .I(data_0)
  ,.C(1'b1)
  ,.IO(o_data[0])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data[2]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB8_D03N")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data_2_iob (
   .I(data_2)
  ,.C(1'b1)
  ,.IO(o_data[2])
);

NX_IOB_O
  // module:~
  // native(1'b0)
  // ring('d0)
  // mandatory(1'b0)
  // protect(1'b0)
  // map_hdlports("IO£o_data1[4]")
  // alias_vhdl("NX_IOB_O")
  // alias_vlog("")
  #(
   .location("IOB9_D01P")
  ,.differential("")
  ,.slewRate("")
  ,.termination("")
  ,.terminationReference("")
  ,.turbo("")
  ,.weakTermination("")
  ,.inputDelayLine("")
  ,.outputDelayLine("")
  ,.inputSignalSlope("")
  ,.outputCapacity("")
  ,.extra('d2)
  ,.locked(1'b0)
  ,.standard("")
  ,.drive("")
  ,.inputDelayOn("")
  ,.outputDelayOn("")
  ,.dynDrive("")
  ,.dynInput("")
  ,.dynTerm("")
  )
  i_o_data1_4_iob (
   .I(data1_4)
  ,.C(1'b1)
  ,.IO(o_data1[4])
);

endmodule
